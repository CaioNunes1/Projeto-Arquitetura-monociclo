// Universidade Federal Rural de Pernambuco
// 2021.2
// Arquitetura e Organização de Computadores - 2ªVA
// Alunos:
// Steffano Pereira
// Haga Fedra
// João Carvalho
// Julyanne Correia
// -----------------------------
`include "i_mem.v"
`include "pc.v"
`include "regfile.v"
`include "ula.v"
`include "sign_extend.v"
`include "d_mem.v"
`include "control/control.v"
`include "jump/jump.v"
`include "utils/utils.v"

module mips(
    input wire clock,
    input wire reset,
    output wire [31:0] nextPC,
    output wire [31:0] ula_result,
    output wire [31:0] data_mem
);

    // ---------------------------------------------
    // Módulo de Controle
    // ---------------------------------------------
    wire MemRead, MemtoReg, MemWrite, ALUSrc, RegWrite, isJAL, isSigned;
    wire [1:0] PCOp, RegDst;

    control mips_control (
        instruction[31:26],
        RegDst,
        PCOp,
        MemRead,
        MemtoReg,
        ula_operation,
        MemWrite,
        ALUSrc,
        RegWrite,
        isJAL,
        isSigned
    );

    // ---------------------------------------------
    // Estágio de Busca de Instruções
    // ---------------------------------------------
    wire [31:0] pc;
    PC pc_check(nextPC, pc, clock);  // Armazena e atualiza o PC

    wire [31:0] pc_increment;  // Representa o valor incrementado do PC
    Adder pc_counter(pc, pc_increment);  // Incrementa o PC

    wire [31:0] instruction;
    i_mem current_instruction(pc, instruction);  // Busca a instrução da memória

    // ---------------------------------------------
    // Estágio de Decodificação
    // ---------------------------------------------
    wire [2:0] ula_operation;
    ula_control mips_ula_control(ula_operation, instruction[5:0], OP);  // Gera sinais de controle da ALU

    // ---------------------------------------------
    // Estágio de Execução
    // ---------------------------------------------
    wire [31:0] ReadData1, ReadData2;
    regfile mips_regfile(
        instruction[25:21],
        instruction[20:16],
        ReadData1,
        ReadData2,
        clock,
        imem_mux_to_write_register,
        to_write_data,
        RegWrite,
        reset
    );  // Lê dados dos registradores

    wire [31:0] regfile_mux_to_ula_In2;
    wire [31:0] sign_extend_to_mux;
    sign_extend mips_sign_extend(instruction[15:0], isSigned, sign_extend_to_mux);  // Extende os valores imediatos com sinal

    mux_32 regfile_mux(ReadData2, sign_extend_to_mux, ALUSrc, regfile_mux_to_ula_In2);  // Seleciona a entrada da ALU

    wire [3:0] OP;
    wire ula_zero_flag;
    ula mips_ula(ReadData1, regfile_mux_to_ula_In2, OP, instruction[10:6], ula_result, ula_zero_flag);  // Executa operações da ALU

    // ---------------------------------------------
    // Estágio de Acesso à Memória
    // ---------------------------------------------
    d_mem mips_d_mem(ula_result, ReadData2, data_mem, MemWrite, MemRead, clock);  // Acessa a memória de dados

    wire [31:0] WriteData;
    mux_32 mux_32_d_mem(ula_result, data_mem, MemtoReg, WriteData);  // Seleciona dados para writeback

    // ---------------------------------------------
    // Estágio de Writeback
    // ---------------------------------------------
    wire [4:0] imem_mux_to_write_register;
    mux_5_4 imem_reg_mux(instruction[20:16], instruction[15:11], 5'b11111, RegDst, imem_mux_to_write_register);

     wire [31:0] to_write_data;
    Adder jal (pc_increment, to_write_data_mux_in2);  // Soma PC para instruções JAL
    mux_32 write_data_mux(WriteData, to_write_data_mux_in2, isJAL, to_write_data);  // Seleciona dados para writeback (JAL ou registrador)

    // ---------------------------------------------
    // Módulo Regfile
    // ---------------------------------------------
    wire [31:0] add_branching_to_mux;
    PCControl pc_control(PCOp, ula_zero_flag, PCSource);  // Gera sinal de controle para o PC baseado em flags e PCOp

    // ---------------------------------------------
    // Módulo de JUMP
    // ---------------------------------------------
    wire [31:0] jump_module_to_mux;
    jump mips_jump(pc_increment[31:28], instruction[25:0], jump_module_to_mux);  // Calcula endereço de salto

    // ---------------------------------------------
    // Módulo de Controle JR
    // ---------------------------------------------
    wire [31:0] jr_PC;
    jr_control mips_jr_control(ula_operation, instruction[5:0], ReadData1, jr_PC);  // Calcula endereço de salto basedado em JR

    // ---------------------------------------------
    // Próximo PC
    // ---------------------------------------------
    wire [1:0] PCSource;  // Sinal de controle para o PC
    mux_32_4 pc_mux (pc_increment, add_branching_to_mux, jump_module_to_mux, jr_PC, PCSource, nextPC);  // Seleciona o próximo PC baseado em vários fatores

endmodule